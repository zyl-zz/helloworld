module test(
	output wire a,
	input wire b
);

assign a = b;

endmodule